BZh91AY&SY��� _�Px��g߰����P{҆0 JB��I�x���i� �z��z���L� �LL&4��!$h�$m@Q�@ ���9�L�����a0CLM0D��M44�2��4  �dh�`{P(������46 m��d��;X^&	��(��:�!�ٵĐ��]~:��`cg[��lf�J���|�4wWn��Y��tl���i�fs}2�I �0߬�^�	�*/+�9,���t�8`	���b�C�j�r\n����f����fXA��l(pZw��Y�\�cN�2s�:���|9HFM��N͊,<�޿/�0J�/�S(߮��D���8�8��41�{�s���(r�K�3�z���܂Ӆ�5��������S��-�nE�H8�z�R�2W�kN0���� t$U,�I�a�P����ҟb������A'�!��g�����6X��$���Jʷ���h��G�<��9��5�F!�)&��1��6ĐTV��u
Ⱥ��K�bq�e֖ad��աPc�XUH��05�e�P1��-�A7��TJ�@3�����\�(�Z���*��O��2�gS��Dt.���$�>&��+�Q�R������d�J'� ���lL�͡Р,�ɋWD
�BrLM�D�y��j%
�aCno�6{�^����+����VaC��8�`;0��elu��iF<�*��abrG�n��3�@�Z#:ٯ[��\m�}�W7J�a�(<�K�һ�<�k2)�\	"9���Q�[���l����t�/4ia���)Q��?��0̃`��E���)����