BZh91AY&SY1y ?_�Py���߰?���P��  �`LM&L�LM2100���&L�20�&�db``9�14L�2da0M4����"RH�@4i�C��  4 D&����ѡ�OMM��i��z�MB5��\Q
 ࣊�兢����?��a�ȠF)��q`��݀`�x�E�T��؊����S=�٣C��W $ b���}'$�˭��t5t�J�nd�_�5(�e�7�{;�������eP7q ��[�O/���7��F��˿��-��tz�����`:!+����6��0p�B0�C ����15��
�%C�d=i�Ļ,�!Q��
�ln~�s`F%>b�:P�d!!$�"a�Iv,_��
Q�	fR��HK��(5��~Vg)����f�
P�BR�6U�	_�fS2�!0�� e	�?�t�Z(<�oe)|>��ߗ,�&~Ad��}��=ߵ>����^5���g����>X�rN� ��A���	��@�Y�7�3���e����T���~X�Z����2�-F�hС�S���n�a=��� }9�#*@� ir*[�|\q`J%��m_��@���0á����l��+X!c�o���N!W�)�(	=��Hj�ˀD�5�ؐi�d���Jd��U�t*��j�x�@؇�]�l�S�y����5}>� �m܄�!x�@w����C�y�!T��/�̗ <
+�@O.�7��lN��7f��x�o �����@���S�p[�|@߬"��=j������5m��KPs�q�4�x�ڍ7A �H0�mA4H*>[GZ Ub��� d!y� YK�X	]�B��T9�h��@\;]}n�P{ (����]�k��'��ɐ���2F�c5�r�[���p	J�AM\�ҁ|$ ��	�~�!�z��Üh����gd��	x=�ttu�pe[�i�5K4�/��j�z�8s�tK���s�@l�6u��@��䔠��t�Ք5l9�HH�����5K^��{d�D�J���b�]��B@X@��